module fa_v2(a,b,ci,s); // fa_v2 module
input a,b,ci; //input
output s; //co가 없음 
wire sm;
_xor2 U0_xor2(.a(a),.b(b),.y(sm));
_xor2 U1_xor2(.a(sm),.b(ci),.y(s));
//instance of xor
endmodule 